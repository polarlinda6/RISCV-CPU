`include "define.v"

module branch_predictor(
	input  clk,
	input  rst_n,
	input  PL_stall,
	input  PL_flush,	
	input  jalr_prediction_en,
	input  B_type_prediction_en,

	output [31:0]jalr_pc_prediction,
	output B_type_prediction_result,

	//jalr
	input  jal,
	input  jalr,
	input  [4:0]Rd,
	input  [31:0]pc_add_4,
	
	input  jal_id,
	input  jalr_id,
	input  [4:0]Rd_id,	
	input  [4:0]Rs1_id,

	//B_type
	input  [31:0]imme,

	input  B_type, 
	input  beq,
	input  bne,
	input  blt,
	input  bge,
	input  bltu,
	input  bgeu,
	input  [31:0]pc,
	input  corrected_result,

	input  B_type_id,
	input  beq_id,
	input  bne_id,
	input  blt_id,
	input  bge_id,
	input  bltu_id,
	input  bgeu_id,
	input  [31:0]pc_id,
	input  B_type_prediction_result_id, 

	input  B_type_branch_failed,
	input  beq_branch_failed,
	input  bne_branch_failed,
	input  blt_branch_failed,
	input  bge_branch_failed,
	input  bltu_branch_failed,
	input  bgeu_branch_failed,
	input  [31:0]pc_branch_filled,
	input  B_type_prediction_result_branch_failed
);

	localparam RAS_STACK_ADDR_WIDTH = 4;

	localparam GHP_INDEX_HR_WIDTH = 6;
	localparam GHP_INDEX_PC_WIDTH = 4;
	localparam LHP_INDEX_HR_WIDTH = 5;
	localparam LHP_INDEX_PC_WIDTH = 3;
	localparam STAT_COUNTER_WIDTH = 4;

	localparam JUMP_STATUS_COUNTER_WIDTH = 2;
	localparam JUMP_STATUS_COUNTER_WIDTH_UB = JUMP_STATUS_COUNTER_WIDTH - 1;


	wire SP_prediction_result;
	wire SP_prediction_result_id;
	wire SP_prediction_result_ex;

	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]GHP_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]GHP_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]GHP_count_ex;

	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_beq_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bne_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_blt_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bge_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bltu_count;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bgeu_count;

	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_beq_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bne_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_blt_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bge_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bltu_count_id;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bgeu_count_id;

	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_beq_count_ex;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bne_count_ex;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_blt_count_ex;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bge_count_ex;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bltu_count_ex;
	wire [JUMP_STATUS_COUNTER_WIDTH_UB:0]LHP_bgeu_count_ex;


	wire GHP_rollback_en_id;
	wire GHP_rollback_en_ex;

	wire GHP_beq_rollback_en_id;
	wire GHP_bne_rollback_en_id;
	wire GHP_blt_rollback_en_id;
	wire GHP_bge_rollback_en_id;
	wire GHP_bltu_rollback_en_id;
	wire GHP_bgeu_rollback_en_id;

	wire GHP_beq_rollback_en_ex;
	wire GHP_bne_rollback_en_ex;
	wire GHP_blt_rollback_en_ex;
	wire GHP_bge_rollback_en_ex;
	wire GHP_bltu_rollback_en_ex;
	wire GHP_bgeu_rollback_en_ex;

	wire LHP_beq_rollback_en_id;
	wire LHP_bne_rollback_en_id;
	wire LHP_blt_rollback_en_id;
	wire LHP_bge_rollback_en_id;
	wire LHP_bltu_rollback_en_id;
	wire LHP_bgeu_rollback_en_id;

	wire LHP_beq_rollback_en_ex;
	wire LHP_bne_rollback_en_ex;
	wire LHP_blt_rollback_en_ex;
	wire LHP_bge_rollback_en_ex;
	wire LHP_bltu_rollback_en_ex;
	wire LHP_bgeu_rollback_en_ex;


	//MP
	meta_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.STAT_COUNTER_WIDTH(STAT_COUNTER_WIDTH)
	) MP_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.prediction_result(B_type_prediction_result),
		.prediction_result_id(B_type_prediction_result_id), 

		.prediction_en(B_type_prediction_en),

		.GHP_beq_rollback_en_id(GHP_beq_rollback_en_id),
		.GHP_bne_rollback_en_id(GHP_bne_rollback_en_id),
		.GHP_blt_rollback_en_id(GHP_blt_rollback_en_id),
		.GHP_bge_rollback_en_id(GHP_bge_rollback_en_id),
		.GHP_bltu_rollback_en_id(GHP_bltu_rollback_en_id),
		.GHP_bgeu_rollback_en_id(GHP_bgeu_rollback_en_id),

		.GHP_beq_rollback_en_ex(GHP_beq_rollback_en_ex),
		.GHP_bne_rollback_en_ex(GHP_bne_rollback_en_ex),
		.GHP_blt_rollback_en_ex(GHP_blt_rollback_en_ex),
		.GHP_bge_rollback_en_ex(GHP_bge_rollback_en_ex),
		.GHP_bltu_rollback_en_ex(GHP_bltu_rollback_en_ex),
		.GHP_bgeu_rollback_en_ex(GHP_bgeu_rollback_en_ex),

		.LHP_beq_rollback_en_id(LHP_beq_rollback_en_id),
		.LHP_bne_rollback_en_id(LHP_bne_rollback_en_id),
		.LHP_blt_rollback_en_id(LHP_blt_rollback_en_id),
		.LHP_bge_rollback_en_id(LHP_bge_rollback_en_id),
		.LHP_bltu_rollback_en_id(LHP_bltu_rollback_en_id),
		.LHP_bgeu_rollback_en_id(LHP_bgeu_rollback_en_id),

		.LHP_beq_rollback_en_ex(LHP_beq_rollback_en_ex),
		.LHP_bne_rollback_en_ex(LHP_bne_rollback_en_ex),
		.LHP_blt_rollback_en_ex(LHP_blt_rollback_en_ex),
		.LHP_bge_rollback_en_ex(LHP_bge_rollback_en_ex),
		.LHP_bltu_rollback_en_ex(LHP_bltu_rollback_en_ex),
		.LHP_bgeu_rollback_en_ex(LHP_bgeu_rollback_en_ex),

		.beq(beq),
		.bne(bne),
		.blt(blt),
		.bge(bge),
		.bltu(bltu),
		.bgeu(bgeu),

		.beq_id(beq_id),  
		.bne_id(bne_id),
		.blt_id(blt_id),
		.bge_id(bge_id),
		.bltu_id(bltu_id),
		.bgeu_id(bgeu_id),

		.beq_ex(beq_ex),
		.bne_ex(bne_ex),
		.blt_ex(blt_ex),
		.bge_ex(bge_ex),
		.bltu_ex(bltu_ex),
		.bgeu_ex(bgeu_ex),

		.SP_prediction_result(SP_prediction_result),
		.SP_prediction_result_id(SP_prediction_result_id),
		.SP_prediction_result_ex(SP_prediction_result_ex),

		.GHP_count(GHP_count),
		.GHP_count_id(GHP_count_id),
		.GHP_count_ex(GHP_count_ex),

		.LHP_beq_count(LHP_beq_count),
		.LHP_bne_count(LHP_bne_count),
		.LHP_blt_count(LHP_blt_count),
		.LHP_bge_count(LHP_bge_count),
		.LHP_bltu_count(LHP_bltu_count),
		.LHP_bgeu_count(LHP_bgeu_count),

		.LHP_beq_count_id(LHP_beq_count_id),
		.LHP_bne_count_id(LHP_bne_count_id),
		.LHP_blt_count_id(LHP_blt_count_id),
		.LHP_bge_count_id(LHP_bge_count_id),
		.LHP_bltu_count_id(LHP_bltu_count_id),
		.LHP_bgeu_count_id(LHP_bgeu_count_id),

		.LHP_beq_count_ex(LHP_beq_count_ex),
		.LHP_bne_count_ex(LHP_bne_count_ex),
		.LHP_blt_count_ex(LHP_blt_count_ex),
		.LHP_bge_count_ex(LHP_bge_count_ex),
		.LHP_bltu_count_ex(LHP_bltu_count_ex),
		.LHP_bgeu_count_ex(LHP_bgeu_count_ex)
	);



	//SP
	static_predictor SP_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.imme_sig(imme[31]),
		.SP_prediction_result(SP_prediction_result),
		.SP_prediction_result_id(SP_prediction_result_id),
		.SP_prediction_result_ex(SP_prediction_result_ex)
	);


	//GHP
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(GHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(GHP_INDEX_PC_WIDTH)
	) GHP_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(B_type),
		.rollback_en_id(GHP_rollback_en_id),
		.rollback_en_ex(GHP_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(GHP_count),
		.HP_count_id(GHP_count_id),
		.HP_count_ex(GHP_count_ex)
	);


	//LHP beq
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_beq_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(beq),
		.rollback_en_id(LHP_beq_rollback_en_id),
		.rollback_en_ex(LHP_beq_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_beq_count),
		.HP_count_id(LHP_beq_count_id),
		.HP_count_ex(LHP_beq_count_ex)
	);
	

	//LHP bne
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_bne_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(bne),
		.rollback_en_id(LHP_bne_rollback_en_id),
		.rollback_en_ex(LHP_bne_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_bne_count),
		.HP_count_id(LHP_bne_count_id),
		.HP_count_ex(LHP_bne_count_ex)
	);
	

	//LHP blt
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_blt_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(blt),
		.rollback_en_id(LHP_blt_rollback_en_id),
		.rollback_en_ex(LHP_blt_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_blt_count),
		.HP_count_id(LHP_blt_count_id),
		.HP_count_ex(LHP_blt_count_ex)
	);
	

	//LHP bge
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_bge_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(bge),
		.rollback_en_id(LHP_bge_rollback_en_id),
		.rollback_en_ex(LHP_bge_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_bge_count),
		.HP_count_id(LHP_bge_count_id),
		.HP_count_ex(LHP_bge_count_ex)
	);
	
	
	//LHP bltu
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_bltu_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(bltu),
		.rollback_en_id(LHP_bltu_rollback_en_id),
		.rollback_en_ex(LHP_bgeu_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_bltu_count),
		.HP_count_id(LHP_bltu_count_id),
		.HP_count_ex(LHP_bltu_count_ex)
	);


	//LHP bgeu
	history_predictor #(
		.JUMP_STATUS_COUNTER_WIDTH(JUMP_STATUS_COUNTER_WIDTH),
		.INDEX_HR_WIDTH(LHP_INDEX_HR_WIDTH),
		.INDEX_PC_WIDTH(LHP_INDEX_PC_WIDTH)
	) LHP_bgeu_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_stall(PL_stall),

		.corrected_result(corrected_result),

		.corrected_en(bgeu),
		.rollback_en_id(LHP_bgeu_rollback_en_id),
		.rollback_en_ex(LHP_bgeu_rollback_en_ex),

		.pc(pc),
		.pc_id(pc_id),
		.pc_ex(pc_branch_filled),

		.HP_count(LHP_bgeu_count),
		.HP_count_id(LHP_bgeu_count_id),
		.HP_count_ex(LHP_bgeu_count_ex)
	);


/////////////////////////////////////////////////////////////////////////////////

	ras #(
		.STACK_ADDR_WIDTH(RAS_STACK_ADDR_WIDTH)
	) ras_inst(
		.clk(clk),
		.rst_n(rst_n),
		.PL_flush(PL_flush),
		.prediction_en(jalr_prediction_en),
		.jal(jal),
		.jalr(jalr),
		.Rd_is_ra(Rd == `ra),
		.pc_add_4(pc_add_4),
		.jal_id(jal_id),
		.jalr_id(jalr_id),
		.Rd_is_ra_id(Rd_id == `ra),
		.Rs1_is_ra_id(Rs1_id == `ra),
		.jalr_pc_prediction(jalr_pc_prediction)
	);

/////////////////////////////////////////////////////////////////////////////////

	wire GHP_failed_en;
	assign GHP_failed_en = B_type_prediction_result_branch_failed == GHP_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB];

	assign GHP_rollback_en_id = PL_flush && B_type_id;
	assign GHP_rollback_en_ex = PL_flush && B_type_branch_failed && GHP_failed_en;

	assign GHP_beq_rollback_en_id  = PL_flush && beq_id;
	assign GHP_bne_rollback_en_id  = PL_flush && bne_ex;
	assign GHP_blt_rollback_en_id  = PL_flush && blt_id;
	assign GHP_bge_rollback_en_id  = PL_flush && bge_id;
	assign GHP_bltu_rollback_en_id = PL_flush && bltu_id;
	assign GHP_bgeu_rollback_en_id = PL_flush && bgeu_id;

	assign GHP_beq_rollback_en_ex  = PL_flush && beq_ex  && GHP_failed_en;
	assign GHP_bne_rollback_en_ex  = PL_flush && bne_ex  && GHP_failed_en;
	assign GHP_blt_rollback_en_ex  = PL_flush && blt_ex  && GHP_failed_en;
	assign GHP_bge_rollback_en_ex  = PL_flush && bge_ex  && GHP_failed_en;
	assign GHP_bltu_rollback_en_ex = PL_flush && bltu_ex && GHP_failed_en;
	assign GHP_bgeu_rollback_en_ex = PL_flush && bgeu_ex && GHP_failed_en;


	assign LHP_beq_rollback_en_id  = PL_flush && beq_id;
	assign LHP_bne_rollback_en_id  = PL_flush && bne_id;
	assign LHP_blt_rollback_en_id  = PL_flush && blt_id;
	assign LHP_bge_rollback_en_id  = PL_flush && bge_id;
	assign LHP_bltu_rollback_en_id = PL_flush && bltu_id;
	assign LHP_bgeu_rollback_en_id = PL_flush && bgeu_id;

	assign LHP_beq_rollback_en_ex  = PL_flush && beq_ex  && (B_type_prediction_result_branch_failed == LHP_beq_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
	assign LHP_bne_rollback_en_ex  = PL_flush && bne_ex  && (B_type_prediction_result_branch_failed == LHP_bne_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
	assign LHP_blt_rollback_en_ex  = PL_flush && blt_ex  && (B_type_prediction_result_branch_failed == LHP_blt_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
	assign LHP_bge_rollback_en_ex  = PL_flush && bge_ex  && (B_type_prediction_result_branch_failed == LHP_bge_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
	assign LHP_bltu_rollback_en_ex = PL_flush && bltu_ex && (B_type_prediction_result_branch_failed == LHP_bltu_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
	assign LHP_bgeu_rollback_en_ex = PL_flush && bgeu_ex && (B_type_prediction_result_branch_failed == LHP_bgeu_count_ex[JUMP_STATUS_COUNTER_CAPACITY_UB]);
endmodule


module static_predictor(
	input clk,
	input rst_n,
	input PL_stall,

	input imme_sig,
	output SP_prediction_result, 
	output SP_prediction_result_id,
	output SP_prediction_result_ex
);
	reg prediciont_result_reg_id, prediciont_result_reg_ex;

	always @(posedge clk)
	begin
		if (!rst_n)
			begin
				prediciont_result_reg_id <= `zero;
				prediciont_result_reg_ex <= `zero;
			end
		else
			begin
				if(!PL_stall)
				begin
					prediciont_result_reg_id <= SP_prediction_result;
					prediciont_result_reg_ex <= prediciont_result_reg_id;
				end
			end
	end	

	assign SP_prediction_result_id = prediciont_result_reg_id;
	assign SP_prediction_result_ex = prediciont_result_reg_ex;
	assign SP_prediction_result = imme_sig;
endmodule